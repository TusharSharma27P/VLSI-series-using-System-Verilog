module AND_GATE(
input a,b,
output y
);
 assign y= a&b;
endmodule
